MIDlet-1: Vocab_en_sv,,br.boirque.vocabuilder.view.Vocabuilder
MIDlet-Data-Size: 51794
MIDlet-Description: Portable Flash Cards to aid on vocabulary learning
MIDlet-Info-URL: http://code.google.com/p/vocabuilder/
MIDlet-Jar-URL: Vocabuilder16_en_sv.jar
MIDlet-Name: Vocabuilder ENGLISH - SWEDISH
MIDlet-Vendor: Cleber Goncalves - Boirque
MIDlet-Version: 1.6.25
MicroEdition-Configuration: CLDC-1.0
MicroEdition-Profile: MIDP-2.0
